module Test(
    input wire clk,
    input wire rst
);

always @(posedge clk) begin
end

endmodule